// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/unisims/STARTUP_FPGACORE.v,v 1.3 2011/05/05 17:01:42 vandanad Exp $
/*

FUNCTION	: Special Function Cell, STARTUP_FPGACORE

*/

`timescale  100 ps / 10 ps

module STARTUP_FPGACORE (CLK, GSR);

    input  CLK, GSR;

endmodule

