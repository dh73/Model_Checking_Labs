// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/unisims/IDELAYCTRL.v,v 1.1 2005/05/10 01:20:05 wloo Exp $

`timescale 1 ps / 1 ps 

module IDELAYCTRL (RDY, REFCLK, RST);

    output RDY;
    input REFCLK;
    input RST;

endmodule // IDELAYCTRL
