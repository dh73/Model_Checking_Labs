// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/unisims/BUFIO.v,v 1.1 2005/05/10 01:20:03 wloo Exp $

`timescale  100 ps / 10 ps

module BUFIO (O, I);

    output O;
    input  I;

endmodule
