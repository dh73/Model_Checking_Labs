// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/unisims/CONFIG.v,v 1.1 2005/05/10 01:20:03 wloo Exp $
`celldefine
`timescale  100 ps / 10 ps

module CONFIG ();

endmodule

