// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/unisims/USR_ACCESS_VIRTEX4.v,v 1.1 2005/05/10 01:20:09 wloo Exp $

`timescale  100 ps / 10 ps

module USR_ACCESS_VIRTEX4 (DATA, DATAVALID);

    output [31:0] DATA;
    output DATAVALID;

endmodule // USR_ACCESS_VIRTEX4
