// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/unisims/CAPTURE_VIRTEX4.v,v 1.1 2005/05/10 01:20:03 wloo Exp $

`timescale  100 ps / 10 ps

module CAPTURE_VIRTEX4 (CAP, CLK);

    input  CAP, CLK;
    parameter ONESHOT = "TRUE";

endmodule
