// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/unisims/STARTUP_SPARTAN3E.v,v 1.1 2005/05/10 01:20:09 wloo Exp $

`timescale  100 ps / 10 ps

module STARTUP_SPARTAN3E (CLK, GSR, GTS, MBT);

    input  CLK, GSR, GTS, MBT;

endmodule
