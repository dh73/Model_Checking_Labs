// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/unisims/FMAP.v,v 1.1 2005/05/10 01:20:03 wloo Exp $

/*

FUNCTION	: FMAP dummy simulation module

*/

`celldefine
`timescale  100 ps / 10 ps

module FMAP (I1, I2, I3, I4, O);

    input  I1, I2, I3, I4, O;

endmodule
