// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/unisims/BUFGMUX_VIRTEX4.v,v 1.1 2005/05/10 01:20:03 wloo Exp $

`timescale 1 ps / 1 ps 

module BUFGMUX_VIRTEX4 (O, I0, I1, S);

    output O;
    input  I0;
    input  I1;
    input  S;

endmodule
