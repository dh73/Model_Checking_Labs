// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/xec_libs/data/unisims/USR_ACCESSE2.v,v 1.1 2010/11/23 20:34:48 vandanad Exp $
///////////////////////////////////////////////////////
//  Copyright (c) 2009 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /     Vendor      : Xilinx 
// \  \    \/      Version     :  12.1
//  \  \           Description : 
//  /  /                      
// /__/   /\       Filename    : Xilinx Formal Library Component - USR_ACCESSE2.v
// \  \  /  \ 
//  \__\/\__ \                    
//                                 
//  Generated by :	/home/chen/xfoundry/HEAD/env/Databases/CAEInterfaces/LibraryWriters/bin/ltw.pl
//  Revision:		1.0
///////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

module USR_ACCESSE2 (
  CFGCLK,
  DATA,
  DATAVALID
);

  output CFGCLK;
  output DATAVALID;
  output [31:0] DATA;


endmodule
